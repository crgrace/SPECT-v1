// File Name: regfile_assign.sv
// Engineer:  Carl Grace (crgrace@lbl.gov)
// Description:  Code used in regfile.sv for assignment
//          
///////////////////////////////////////////////////////////////////

config_bits[BYPASS_SEL] <= 8'h00;
config_bits[EXT_RESET_0] <= 8'h00;
config_bits[EXT_RESET_1] <= 8'h00;
config_bits[EXT_RESET_2] <= 8'h00;
config_bits[FB_DEL_CTRL] <= 8'hFF;
config_bits[GAIN_SEL] <= 8'h00;
config_bits[PD_ANODE_0] <= 8'h00;
config_bits[PD_ANODE_1] <= 8'h00;
config_bits[PD_CATHODE_RST_SEL] <= 8'h00;


